module IDEX(
    CLK,
    
)