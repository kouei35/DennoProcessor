module EXMEM(

);