module test_IDEX();

