module rs1mux(
    rs1muxsel,
    rs1val,
    ALUOUT,
    PC
);

