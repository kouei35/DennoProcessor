module FowardingAdjustUnit2(

);