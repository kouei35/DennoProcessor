module EXMEM(
    ALUOUT,
    Z_flag,
    PC,
    DmemREB,
    DmemWEB,
    
);