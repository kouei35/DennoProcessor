module IDEX_test();

ControlUnit ControlUnit();
regfile regfile();
LoadStoremux LoadStoremux();
twelve2thirtytwosext twelve2thirtytwosext();
twenty2thirtytwosext twenty2thirtytwosext();
mux2 mux2();
shifer1 shifer1();
shifer12 shifer12();
IDEX IDEX();

IFIDBlock IFIDBlock();